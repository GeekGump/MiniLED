module gw_gao(
    app_en,
    \app_cmd[2] ,
    \app_cmd[1] ,
    \app_cmd[0] ,
    \app_addr[27] ,
    \app_addr[26] ,
    \app_addr[25] ,
    \app_addr[24] ,
    \app_addr[23] ,
    \app_addr[22] ,
    \app_addr[21] ,
    \app_addr[20] ,
    \app_addr[19] ,
    \app_addr[18] ,
    \app_addr[17] ,
    \app_addr[16] ,
    \app_addr[15] ,
    \app_addr[14] ,
    \app_addr[13] ,
    \app_addr[12] ,
    \app_addr[11] ,
    \app_addr[10] ,
    \app_addr[9] ,
    \app_addr[8] ,
    \app_addr[7] ,
    \app_addr[6] ,
    \app_addr[5] ,
    \app_addr[4] ,
    \app_addr[3] ,
    \app_addr[2] ,
    \app_addr[1] ,
    \app_addr[0] ,
    app_wdf_rdy,
    app_rdy,
    app_wdf_wren,
    app_wdf_end,
    \app_wdf_data[63] ,
    \app_wdf_data[62] ,
    \app_wdf_data[61] ,
    \app_wdf_data[60] ,
    \app_wdf_data[59] ,
    \app_wdf_data[58] ,
    \app_wdf_data[57] ,
    \app_wdf_data[56] ,
    \app_wdf_data[55] ,
    \app_wdf_data[54] ,
    \app_wdf_data[53] ,
    \app_wdf_data[52] ,
    \app_wdf_data[51] ,
    \app_wdf_data[50] ,
    \app_wdf_data[49] ,
    \app_wdf_data[48] ,
    \app_wdf_data[47] ,
    \app_wdf_data[46] ,
    \app_wdf_data[45] ,
    \app_wdf_data[44] ,
    \app_wdf_data[43] ,
    \app_wdf_data[42] ,
    \app_wdf_data[41] ,
    \app_wdf_data[40] ,
    \app_wdf_data[39] ,
    \app_wdf_data[38] ,
    \app_wdf_data[37] ,
    \app_wdf_data[36] ,
    \app_wdf_data[35] ,
    \app_wdf_data[34] ,
    \app_wdf_data[33] ,
    \app_wdf_data[32] ,
    \app_wdf_data[31] ,
    \app_wdf_data[30] ,
    \app_wdf_data[29] ,
    \app_wdf_data[28] ,
    \app_wdf_data[27] ,
    \app_wdf_data[26] ,
    \app_wdf_data[25] ,
    \app_wdf_data[24] ,
    \app_wdf_data[23] ,
    \app_wdf_data[22] ,
    \app_wdf_data[21] ,
    \app_wdf_data[20] ,
    \app_wdf_data[19] ,
    \app_wdf_data[18] ,
    \app_wdf_data[17] ,
    \app_wdf_data[16] ,
    \app_wdf_data[15] ,
    \app_wdf_data[14] ,
    \app_wdf_data[13] ,
    \app_wdf_data[12] ,
    \app_wdf_data[11] ,
    \app_wdf_data[10] ,
    \app_wdf_data[9] ,
    \app_wdf_data[8] ,
    \app_wdf_data[7] ,
    \app_wdf_data[6] ,
    \app_wdf_data[5] ,
    \app_wdf_data[4] ,
    \app_wdf_data[3] ,
    \app_wdf_data[2] ,
    \app_wdf_data[1] ,
    \app_wdf_data[0] ,
    app_rd_data_valid,
    app_rd_data_end,
    \app_rd_data[63] ,
    \app_rd_data[62] ,
    \app_rd_data[61] ,
    \app_rd_data[60] ,
    \app_rd_data[59] ,
    \app_rd_data[58] ,
    \app_rd_data[57] ,
    \app_rd_data[56] ,
    \app_rd_data[55] ,
    \app_rd_data[54] ,
    \app_rd_data[53] ,
    \app_rd_data[52] ,
    \app_rd_data[51] ,
    \app_rd_data[50] ,
    \app_rd_data[49] ,
    \app_rd_data[48] ,
    \app_rd_data[47] ,
    \app_rd_data[46] ,
    \app_rd_data[45] ,
    \app_rd_data[44] ,
    \app_rd_data[43] ,
    \app_rd_data[42] ,
    \app_rd_data[41] ,
    \app_rd_data[40] ,
    \app_rd_data[39] ,
    \app_rd_data[38] ,
    \app_rd_data[37] ,
    \app_rd_data[36] ,
    \app_rd_data[35] ,
    \app_rd_data[34] ,
    \app_rd_data[33] ,
    \app_rd_data[32] ,
    \app_rd_data[31] ,
    \app_rd_data[30] ,
    \app_rd_data[29] ,
    \app_rd_data[28] ,
    \app_rd_data[27] ,
    \app_rd_data[26] ,
    \app_rd_data[25] ,
    \app_rd_data[24] ,
    \app_rd_data[23] ,
    \app_rd_data[22] ,
    \app_rd_data[21] ,
    \app_rd_data[20] ,
    \app_rd_data[19] ,
    \app_rd_data[18] ,
    \app_rd_data[17] ,
    \app_rd_data[16] ,
    \app_rd_data[15] ,
    \app_rd_data[14] ,
    \app_rd_data[13] ,
    \app_rd_data[12] ,
    \app_rd_data[11] ,
    \app_rd_data[10] ,
    \app_rd_data[9] ,
    \app_rd_data[8] ,
    \app_rd_data[7] ,
    \app_rd_data[6] ,
    \app_rd_data[5] ,
    \app_rd_data[4] ,
    \app_rd_data[3] ,
    \app_rd_data[2] ,
    \app_rd_data[1] ,
    \app_rd_data[0] ,
    error,
    error_flag,
    \lvds_video_top_inst/max[7] ,
    \lvds_video_top_inst/max[6] ,
    \lvds_video_top_inst/max[5] ,
    \lvds_video_top_inst/max[4] ,
    \lvds_video_top_inst/max[3] ,
    \lvds_video_top_inst/max[2] ,
    \lvds_video_top_inst/max[1] ,
    \lvds_video_top_inst/max[0] ,
    clk_x1,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input app_en;
input \app_cmd[2] ;
input \app_cmd[1] ;
input \app_cmd[0] ;
input \app_addr[27] ;
input \app_addr[26] ;
input \app_addr[25] ;
input \app_addr[24] ;
input \app_addr[23] ;
input \app_addr[22] ;
input \app_addr[21] ;
input \app_addr[20] ;
input \app_addr[19] ;
input \app_addr[18] ;
input \app_addr[17] ;
input \app_addr[16] ;
input \app_addr[15] ;
input \app_addr[14] ;
input \app_addr[13] ;
input \app_addr[12] ;
input \app_addr[11] ;
input \app_addr[10] ;
input \app_addr[9] ;
input \app_addr[8] ;
input \app_addr[7] ;
input \app_addr[6] ;
input \app_addr[5] ;
input \app_addr[4] ;
input \app_addr[3] ;
input \app_addr[2] ;
input \app_addr[1] ;
input \app_addr[0] ;
input app_wdf_rdy;
input app_rdy;
input app_wdf_wren;
input app_wdf_end;
input \app_wdf_data[63] ;
input \app_wdf_data[62] ;
input \app_wdf_data[61] ;
input \app_wdf_data[60] ;
input \app_wdf_data[59] ;
input \app_wdf_data[58] ;
input \app_wdf_data[57] ;
input \app_wdf_data[56] ;
input \app_wdf_data[55] ;
input \app_wdf_data[54] ;
input \app_wdf_data[53] ;
input \app_wdf_data[52] ;
input \app_wdf_data[51] ;
input \app_wdf_data[50] ;
input \app_wdf_data[49] ;
input \app_wdf_data[48] ;
input \app_wdf_data[47] ;
input \app_wdf_data[46] ;
input \app_wdf_data[45] ;
input \app_wdf_data[44] ;
input \app_wdf_data[43] ;
input \app_wdf_data[42] ;
input \app_wdf_data[41] ;
input \app_wdf_data[40] ;
input \app_wdf_data[39] ;
input \app_wdf_data[38] ;
input \app_wdf_data[37] ;
input \app_wdf_data[36] ;
input \app_wdf_data[35] ;
input \app_wdf_data[34] ;
input \app_wdf_data[33] ;
input \app_wdf_data[32] ;
input \app_wdf_data[31] ;
input \app_wdf_data[30] ;
input \app_wdf_data[29] ;
input \app_wdf_data[28] ;
input \app_wdf_data[27] ;
input \app_wdf_data[26] ;
input \app_wdf_data[25] ;
input \app_wdf_data[24] ;
input \app_wdf_data[23] ;
input \app_wdf_data[22] ;
input \app_wdf_data[21] ;
input \app_wdf_data[20] ;
input \app_wdf_data[19] ;
input \app_wdf_data[18] ;
input \app_wdf_data[17] ;
input \app_wdf_data[16] ;
input \app_wdf_data[15] ;
input \app_wdf_data[14] ;
input \app_wdf_data[13] ;
input \app_wdf_data[12] ;
input \app_wdf_data[11] ;
input \app_wdf_data[10] ;
input \app_wdf_data[9] ;
input \app_wdf_data[8] ;
input \app_wdf_data[7] ;
input \app_wdf_data[6] ;
input \app_wdf_data[5] ;
input \app_wdf_data[4] ;
input \app_wdf_data[3] ;
input \app_wdf_data[2] ;
input \app_wdf_data[1] ;
input \app_wdf_data[0] ;
input app_rd_data_valid;
input app_rd_data_end;
input \app_rd_data[63] ;
input \app_rd_data[62] ;
input \app_rd_data[61] ;
input \app_rd_data[60] ;
input \app_rd_data[59] ;
input \app_rd_data[58] ;
input \app_rd_data[57] ;
input \app_rd_data[56] ;
input \app_rd_data[55] ;
input \app_rd_data[54] ;
input \app_rd_data[53] ;
input \app_rd_data[52] ;
input \app_rd_data[51] ;
input \app_rd_data[50] ;
input \app_rd_data[49] ;
input \app_rd_data[48] ;
input \app_rd_data[47] ;
input \app_rd_data[46] ;
input \app_rd_data[45] ;
input \app_rd_data[44] ;
input \app_rd_data[43] ;
input \app_rd_data[42] ;
input \app_rd_data[41] ;
input \app_rd_data[40] ;
input \app_rd_data[39] ;
input \app_rd_data[38] ;
input \app_rd_data[37] ;
input \app_rd_data[36] ;
input \app_rd_data[35] ;
input \app_rd_data[34] ;
input \app_rd_data[33] ;
input \app_rd_data[32] ;
input \app_rd_data[31] ;
input \app_rd_data[30] ;
input \app_rd_data[29] ;
input \app_rd_data[28] ;
input \app_rd_data[27] ;
input \app_rd_data[26] ;
input \app_rd_data[25] ;
input \app_rd_data[24] ;
input \app_rd_data[23] ;
input \app_rd_data[22] ;
input \app_rd_data[21] ;
input \app_rd_data[20] ;
input \app_rd_data[19] ;
input \app_rd_data[18] ;
input \app_rd_data[17] ;
input \app_rd_data[16] ;
input \app_rd_data[15] ;
input \app_rd_data[14] ;
input \app_rd_data[13] ;
input \app_rd_data[12] ;
input \app_rd_data[11] ;
input \app_rd_data[10] ;
input \app_rd_data[9] ;
input \app_rd_data[8] ;
input \app_rd_data[7] ;
input \app_rd_data[6] ;
input \app_rd_data[5] ;
input \app_rd_data[4] ;
input \app_rd_data[3] ;
input \app_rd_data[2] ;
input \app_rd_data[1] ;
input \app_rd_data[0] ;
input error;
input error_flag;
input \lvds_video_top_inst/max[7] ;
input \lvds_video_top_inst/max[6] ;
input \lvds_video_top_inst/max[5] ;
input \lvds_video_top_inst/max[4] ;
input \lvds_video_top_inst/max[3] ;
input \lvds_video_top_inst/max[2] ;
input \lvds_video_top_inst/max[1] ;
input \lvds_video_top_inst/max[0] ;
input clk_x1;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire app_en;
wire \app_cmd[2] ;
wire \app_cmd[1] ;
wire \app_cmd[0] ;
wire \app_addr[27] ;
wire \app_addr[26] ;
wire \app_addr[25] ;
wire \app_addr[24] ;
wire \app_addr[23] ;
wire \app_addr[22] ;
wire \app_addr[21] ;
wire \app_addr[20] ;
wire \app_addr[19] ;
wire \app_addr[18] ;
wire \app_addr[17] ;
wire \app_addr[16] ;
wire \app_addr[15] ;
wire \app_addr[14] ;
wire \app_addr[13] ;
wire \app_addr[12] ;
wire \app_addr[11] ;
wire \app_addr[10] ;
wire \app_addr[9] ;
wire \app_addr[8] ;
wire \app_addr[7] ;
wire \app_addr[6] ;
wire \app_addr[5] ;
wire \app_addr[4] ;
wire \app_addr[3] ;
wire \app_addr[2] ;
wire \app_addr[1] ;
wire \app_addr[0] ;
wire app_wdf_rdy;
wire app_rdy;
wire app_wdf_wren;
wire app_wdf_end;
wire \app_wdf_data[63] ;
wire \app_wdf_data[62] ;
wire \app_wdf_data[61] ;
wire \app_wdf_data[60] ;
wire \app_wdf_data[59] ;
wire \app_wdf_data[58] ;
wire \app_wdf_data[57] ;
wire \app_wdf_data[56] ;
wire \app_wdf_data[55] ;
wire \app_wdf_data[54] ;
wire \app_wdf_data[53] ;
wire \app_wdf_data[52] ;
wire \app_wdf_data[51] ;
wire \app_wdf_data[50] ;
wire \app_wdf_data[49] ;
wire \app_wdf_data[48] ;
wire \app_wdf_data[47] ;
wire \app_wdf_data[46] ;
wire \app_wdf_data[45] ;
wire \app_wdf_data[44] ;
wire \app_wdf_data[43] ;
wire \app_wdf_data[42] ;
wire \app_wdf_data[41] ;
wire \app_wdf_data[40] ;
wire \app_wdf_data[39] ;
wire \app_wdf_data[38] ;
wire \app_wdf_data[37] ;
wire \app_wdf_data[36] ;
wire \app_wdf_data[35] ;
wire \app_wdf_data[34] ;
wire \app_wdf_data[33] ;
wire \app_wdf_data[32] ;
wire \app_wdf_data[31] ;
wire \app_wdf_data[30] ;
wire \app_wdf_data[29] ;
wire \app_wdf_data[28] ;
wire \app_wdf_data[27] ;
wire \app_wdf_data[26] ;
wire \app_wdf_data[25] ;
wire \app_wdf_data[24] ;
wire \app_wdf_data[23] ;
wire \app_wdf_data[22] ;
wire \app_wdf_data[21] ;
wire \app_wdf_data[20] ;
wire \app_wdf_data[19] ;
wire \app_wdf_data[18] ;
wire \app_wdf_data[17] ;
wire \app_wdf_data[16] ;
wire \app_wdf_data[15] ;
wire \app_wdf_data[14] ;
wire \app_wdf_data[13] ;
wire \app_wdf_data[12] ;
wire \app_wdf_data[11] ;
wire \app_wdf_data[10] ;
wire \app_wdf_data[9] ;
wire \app_wdf_data[8] ;
wire \app_wdf_data[7] ;
wire \app_wdf_data[6] ;
wire \app_wdf_data[5] ;
wire \app_wdf_data[4] ;
wire \app_wdf_data[3] ;
wire \app_wdf_data[2] ;
wire \app_wdf_data[1] ;
wire \app_wdf_data[0] ;
wire app_rd_data_valid;
wire app_rd_data_end;
wire \app_rd_data[63] ;
wire \app_rd_data[62] ;
wire \app_rd_data[61] ;
wire \app_rd_data[60] ;
wire \app_rd_data[59] ;
wire \app_rd_data[58] ;
wire \app_rd_data[57] ;
wire \app_rd_data[56] ;
wire \app_rd_data[55] ;
wire \app_rd_data[54] ;
wire \app_rd_data[53] ;
wire \app_rd_data[52] ;
wire \app_rd_data[51] ;
wire \app_rd_data[50] ;
wire \app_rd_data[49] ;
wire \app_rd_data[48] ;
wire \app_rd_data[47] ;
wire \app_rd_data[46] ;
wire \app_rd_data[45] ;
wire \app_rd_data[44] ;
wire \app_rd_data[43] ;
wire \app_rd_data[42] ;
wire \app_rd_data[41] ;
wire \app_rd_data[40] ;
wire \app_rd_data[39] ;
wire \app_rd_data[38] ;
wire \app_rd_data[37] ;
wire \app_rd_data[36] ;
wire \app_rd_data[35] ;
wire \app_rd_data[34] ;
wire \app_rd_data[33] ;
wire \app_rd_data[32] ;
wire \app_rd_data[31] ;
wire \app_rd_data[30] ;
wire \app_rd_data[29] ;
wire \app_rd_data[28] ;
wire \app_rd_data[27] ;
wire \app_rd_data[26] ;
wire \app_rd_data[25] ;
wire \app_rd_data[24] ;
wire \app_rd_data[23] ;
wire \app_rd_data[22] ;
wire \app_rd_data[21] ;
wire \app_rd_data[20] ;
wire \app_rd_data[19] ;
wire \app_rd_data[18] ;
wire \app_rd_data[17] ;
wire \app_rd_data[16] ;
wire \app_rd_data[15] ;
wire \app_rd_data[14] ;
wire \app_rd_data[13] ;
wire \app_rd_data[12] ;
wire \app_rd_data[11] ;
wire \app_rd_data[10] ;
wire \app_rd_data[9] ;
wire \app_rd_data[8] ;
wire \app_rd_data[7] ;
wire \app_rd_data[6] ;
wire \app_rd_data[5] ;
wire \app_rd_data[4] ;
wire \app_rd_data[3] ;
wire \app_rd_data[2] ;
wire \app_rd_data[1] ;
wire \app_rd_data[0] ;
wire error;
wire error_flag;
wire \lvds_video_top_inst/max[7] ;
wire \lvds_video_top_inst/max[6] ;
wire \lvds_video_top_inst/max[5] ;
wire \lvds_video_top_inst/max[4] ;
wire \lvds_video_top_inst/max[3] ;
wire \lvds_video_top_inst/max[2] ;
wire \lvds_video_top_inst/max[1] ;
wire \lvds_video_top_inst/max[0] ;
wire clk_x1;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({app_rd_data_valid,error,error_flag}),
    .trig1_i({\lvds_video_top_inst/max[7] ,\lvds_video_top_inst/max[6] ,\lvds_video_top_inst/max[5] ,\lvds_video_top_inst/max[4] ,\lvds_video_top_inst/max[3] ,\lvds_video_top_inst/max[2] ,\lvds_video_top_inst/max[1] ,\lvds_video_top_inst/max[0] }),
    .data_i({app_en,\app_cmd[2] ,\app_cmd[1] ,\app_cmd[0] ,\app_addr[27] ,\app_addr[26] ,\app_addr[25] ,\app_addr[24] ,\app_addr[23] ,\app_addr[22] ,\app_addr[21] ,\app_addr[20] ,\app_addr[19] ,\app_addr[18] ,\app_addr[17] ,\app_addr[16] ,\app_addr[15] ,\app_addr[14] ,\app_addr[13] ,\app_addr[12] ,\app_addr[11] ,\app_addr[10] ,\app_addr[9] ,\app_addr[8] ,\app_addr[7] ,\app_addr[6] ,\app_addr[5] ,\app_addr[4] ,\app_addr[3] ,\app_addr[2] ,\app_addr[1] ,\app_addr[0] ,app_wdf_rdy,app_rdy,app_wdf_wren,app_wdf_end,\app_wdf_data[63] ,\app_wdf_data[62] ,\app_wdf_data[61] ,\app_wdf_data[60] ,\app_wdf_data[59] ,\app_wdf_data[58] ,\app_wdf_data[57] ,\app_wdf_data[56] ,\app_wdf_data[55] ,\app_wdf_data[54] ,\app_wdf_data[53] ,\app_wdf_data[52] ,\app_wdf_data[51] ,\app_wdf_data[50] ,\app_wdf_data[49] ,\app_wdf_data[48] ,\app_wdf_data[47] ,\app_wdf_data[46] ,\app_wdf_data[45] ,\app_wdf_data[44] ,\app_wdf_data[43] ,\app_wdf_data[42] ,\app_wdf_data[41] ,\app_wdf_data[40] ,\app_wdf_data[39] ,\app_wdf_data[38] ,\app_wdf_data[37] ,\app_wdf_data[36] ,\app_wdf_data[35] ,\app_wdf_data[34] ,\app_wdf_data[33] ,\app_wdf_data[32] ,\app_wdf_data[31] ,\app_wdf_data[30] ,\app_wdf_data[29] ,\app_wdf_data[28] ,\app_wdf_data[27] ,\app_wdf_data[26] ,\app_wdf_data[25] ,\app_wdf_data[24] ,\app_wdf_data[23] ,\app_wdf_data[22] ,\app_wdf_data[21] ,\app_wdf_data[20] ,\app_wdf_data[19] ,\app_wdf_data[18] ,\app_wdf_data[17] ,\app_wdf_data[16] ,\app_wdf_data[15] ,\app_wdf_data[14] ,\app_wdf_data[13] ,\app_wdf_data[12] ,\app_wdf_data[11] ,\app_wdf_data[10] ,\app_wdf_data[9] ,\app_wdf_data[8] ,\app_wdf_data[7] ,\app_wdf_data[6] ,\app_wdf_data[5] ,\app_wdf_data[4] ,\app_wdf_data[3] ,\app_wdf_data[2] ,\app_wdf_data[1] ,\app_wdf_data[0] ,app_rd_data_valid,app_rd_data_end,\app_rd_data[63] ,\app_rd_data[62] ,\app_rd_data[61] ,\app_rd_data[60] ,\app_rd_data[59] ,\app_rd_data[58] ,\app_rd_data[57] ,\app_rd_data[56] ,\app_rd_data[55] ,\app_rd_data[54] ,\app_rd_data[53] ,\app_rd_data[52] ,\app_rd_data[51] ,\app_rd_data[50] ,\app_rd_data[49] ,\app_rd_data[48] ,\app_rd_data[47] ,\app_rd_data[46] ,\app_rd_data[45] ,\app_rd_data[44] ,\app_rd_data[43] ,\app_rd_data[42] ,\app_rd_data[41] ,\app_rd_data[40] ,\app_rd_data[39] ,\app_rd_data[38] ,\app_rd_data[37] ,\app_rd_data[36] ,\app_rd_data[35] ,\app_rd_data[34] ,\app_rd_data[33] ,\app_rd_data[32] ,\app_rd_data[31] ,\app_rd_data[30] ,\app_rd_data[29] ,\app_rd_data[28] ,\app_rd_data[27] ,\app_rd_data[26] ,\app_rd_data[25] ,\app_rd_data[24] ,\app_rd_data[23] ,\app_rd_data[22] ,\app_rd_data[21] ,\app_rd_data[20] ,\app_rd_data[19] ,\app_rd_data[18] ,\app_rd_data[17] ,\app_rd_data[16] ,\app_rd_data[15] ,\app_rd_data[14] ,\app_rd_data[13] ,\app_rd_data[12] ,\app_rd_data[11] ,\app_rd_data[10] ,\app_rd_data[9] ,\app_rd_data[8] ,\app_rd_data[7] ,\app_rd_data[6] ,\app_rd_data[5] ,\app_rd_data[4] ,\app_rd_data[3] ,\app_rd_data[2] ,\app_rd_data[1] ,\app_rd_data[0] ,error,error_flag}),
    .clk_i(clk_x1)
);

endmodule
