//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.03 (64-bit)
//Part Number: GW2A-LV55PG484C8/I7
//Device: GW2A-55
//Device Version: C
//Created Time: Tue Jun 18 16:00:04 2024

module SPI7001_25M_1M_rPLL (clkout, clkoutd, clkin);

output clkout;
output clkoutd;
input clkin;

wire lock_o;
wire clkoutp_o;
wire clkoutd3_o;
wire gw_gnd;

assign gw_gnd = 1'b0;

rPLL  led_rpll_inst(
    .CLKOUT(clkout),
    .LOCK(lock_o),
    .CLKOUTP(clkoutp_o),
    .CLKOUTD(clkoutd),
    .CLKOUTD3(clkoutd3_o),
    .RESET(gw_gnd),
    .RESET_P(gw_gnd),
    .CLKIN(clkin),
    .CLKFB(gw_gnd),
    .FBDSEL({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
    .IDSEL({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
    .ODSEL({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
    .PSDA({gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
    .DUTYDA({gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
    .FDLY({gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam led_rpll_inst.FCLKIN = "50";
defparam led_rpll_inst.DYN_IDIV_SEL = "false";
defparam led_rpll_inst.IDIV_SEL = 1;
defparam led_rpll_inst.DYN_FBDIV_SEL = "false";
defparam led_rpll_inst.FBDIV_SEL = 0;
defparam led_rpll_inst.DYN_ODIV_SEL = "false";
defparam led_rpll_inst.ODIV_SEL = 32;
defparam led_rpll_inst.PSDA_SEL = "0000";
defparam led_rpll_inst.DYN_DA_EN = "true";
defparam led_rpll_inst.DUTYDA_SEL = "1000";
defparam led_rpll_inst.CLKOUT_FT_DIR = 1'b1;
defparam led_rpll_inst.CLKOUTP_FT_DIR = 1'b1;
defparam led_rpll_inst.CLKOUT_DLY_STEP = 0;
defparam led_rpll_inst.CLKOUTP_DLY_STEP = 0;
defparam led_rpll_inst.CLKFB_SEL = "internal";
defparam led_rpll_inst.CLKOUT_BYPASS = "false";
defparam led_rpll_inst.CLKOUTP_BYPASS = "false";
defparam led_rpll_inst.CLKOUTD_BYPASS = "false";
defparam led_rpll_inst.DYN_SDIV_SEL = 26;
defparam led_rpll_inst.CLKOUTD_SRC = "CLKOUT";
defparam led_rpll_inst.CLKOUTD3_SRC = "CLKOUT";
defparam led_rpll_inst.DEVICE = "GW2A-55C";

endmodule //SPI7001_25M_1M_rPLL
